module clk_div_v1 (

);

    always @(posedge sys_clk) begin
        
    end
endmodule