library verilog;
use verilog.vl_types.all;
entity risc_tb is
end risc_tb;
