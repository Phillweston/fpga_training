
module my_issp (
	source,
	probe);	

	output	[10:0]	source;
	input	[0:0]	probe;
endmodule
