library verilog;
use verilog.vl_types.all;
entity digital_clock_v1_tb is
end digital_clock_v1_tb;
