module alu (
    // ????
    input           clk,        // RISC??????
    input           rst_n,      // RISC????????
    // ????????
    input           en_alu,     // en_alu==1??out_alu??
    // ?????
    input [15:13]   ir,         // ?????
    // ??????????
    input [7:0]     bus_data,   // RISC????
    input [7:0]     out_acc,    // ??????
    // ALU??
    output reg [7:0] out_alu    // ALU???
);

	localparam
		// ?????
		NOP     = 3'b000,    // ???
		LDA     = 3'b001,    // ???????????????
		STO     = 3'b010,    // ???????????????
		ADD     = 3'b011,    // ???????????????
		NXOR    = 3'b100,    // ????????????????????
		SFT     = 3'b101,    // ????????????????
		SKP     = 3'b110,    // ???????????????
		NJMP    = 3'b111;    // ????????????

	always @(posedge clk or negedge rst_n) begin
		if (~rst_n)
			out_alu <= 8'd0;
		else if (en_alu)
			case (ir[15:13])
				NOP  : out_alu <= out_alu;
				LDA  : out_alu <= bus_data;
				STO  : out_alu <= out_alu;
				ADD  : out_alu <= bus_data + out_acc;
				NXOR : out_alu <= bus_data ^ out_acc;
				SFT  : out_alu <= {bus_data[6:0], bus_data[7]};
				SKP  : out_alu <= out_alu;
				NJMP : out_alu <= out_alu;
				default : out_alu <= out_alu;
			endcase
	end

endmodule