module led_driver_v3 (

);
reg [31:0] cnt;
endmodule