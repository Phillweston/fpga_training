library verilog;
use verilog.vl_types.all;
entity tesebench is
end tesebench;
