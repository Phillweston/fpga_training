library verilog;
use verilog.vl_types.all;
entity m_seq_gen_test is
end m_seq_gen_test;
