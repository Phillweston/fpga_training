module img_filter
(
	//邻域像素点
	input [7:0]			p00,	//邻域1*1像素点
	input [7:0]			p01,	//邻域1*2像素点
	input [7:0]			p02,	//邻域1*3像素点
	input [7:0]			p10,	//领域2*1像素点
	input [7:0]			p11,	//领域2*2像素点，中心像素点
	input [7:0]			p12,	//领域2*3像素点
	input [7:0]			p20,	//领域3*1像素点
	input [7:0]			p21,	//领域3*2像素点
	input [7:0]			p22,	//领域3*3像素点
	//输出平均值
	output [7:0]		oval	//邻域平均值
);
	//////////////////数学平均/////////////////////////////////////////////////////////
	/*
	wire [11:0]	sum;
	assign sum = p00 + p01 + p02 +
				 p10 + p11 + p12 +
				 p20 + p21 + p22;

	wire [11:0]	oval_r;
	assign oval_r = sum/12'd9;
	assign oval = oval_r[7:0]; */


	//////////////////加权平均//////////////////////////////////////////////////////////////////
	/*
	P00	P01	P02       1	2	1
	P10	P11	P12       2	4	2
	P20	P21	P22       1	2	1
	*/
	/*
	wire [11:0] sub;
	assign sub = ({4'd0,p00[7:0]}<<0) + ({4'd0,p01[7:0]}<<1) + ({4'd0,p02[7:0]}<<0) +
				 ({4'd0,p10[7:0]}<<1) + ({4'd0,p11[7:0]}<<2) + ({4'd0,p12[7:0]}<<1) +
				 ({4'd0,p20[7:0]}<<0) + ({4'd0,p21[7:0]}<<1) + ({4'd0,p22[7:0]}<<0);   
	assign oval = sub[11:4];
	*/

	//第1次遍历/////////////
	wire [7:0] max00,max01,max02,max03,max04,max05,max06,max07;
	wire [7:0] min00,min01,min02,min03,min04,min05,min06,min07;

	switch switch00
	(
		//被比较交换的数输入
		.d0(p00),		//参与交互的第1个数
		.d1(p01),		//参与交互的第2个数
		//输出交互后的数据
		.max(max00),	//交互比较后的最大的数据
		.min(min00)		//交互比较后的最小的数据
	);
	switch switch01
	(
		//被比较交换的数输入
		.d0(max00),		//参与交互的第1个数
		.d1(p02),		//参与交互的第2个数
		//输出交互后的数据
		.max(max01),	//交互比较后的最大的数据
		.min(min01)		//交互比较后的最小的数据
	);
	switch switch02
	(
		//被比较交换的数输入
		.d0(max01),		//参与交互的第1个数
		.d1(p10),		//参与交互的第2个数
		//输出交互后的数据
		.max(max02),	//交互比较后的最大的数据
		.min(min02)		//交互比较后的最小的数据
	);
	switch switch03
	(
		//被比较交换的数输入
		.d0(max02),		//参与交互的第1个数
		.d1(p11),		//参与交互的第2个数
		//输出交互后的数据
		.max(max03),	//交互比较后的最大的数据
		.min(min03)		//交互比较后的最小的数据
	);
	switch switch04
	(
		//被比较交换的数输入
		.d0(max03),		//参与交互的第1个数
		.d1(p12),		//参与交互的第2个数
		//输出交互后的数据
		.max(max04),	//交互比较后的最大的数据
		.min(min04)		//交互比较后的最小的数据
	);
	switch switch05
	(
		//被比较交换的数输入
		.d0(max04),		//参与交互的第1个数
		.d1(p20),		//参与交互的第2个数
		//输出交互后的数据
		.max(max05),	//交互比较后的最大的数据
		.min(min05)		//交互比较后的最小的数据
	);
	switch switch06
	(
		//被比较交换的数输入
		.d0(max05),		//参与交互的第1个数
		.d1(p21),		//参与交互的第2个数
		//输出交互后的数据
		.max(max06),	//交互比较后的最大的数据
		.min(min06)		//交互比较后的最小的数据
	);
	switch switch07
	(
		//被比较交换的数输入
		.d0(max06),		//参与交互的第1个数
		.d1(p22),		//参与交互的第2个数
		//输出交互后的数据
		.max(max07),	//交互比较后的最大的数据
		.min(min07)		//交互比较后的最小的数据
	);

	//第2次遍历/////////////
	wire [7:0] max10,max11,max12,max13,max14,max15,max16;
	wire [7:0] min10,min11,min12,min13,min14,min15,min16;

	switch switch10
	(
		//被比较交换的数输入
		.d0(min00),		//参与交互的第1个数
		.d1(min01),		//参与交互的第2个数
		//输出交互后的数据
		.max(max10),	//交互比较后的最大的数据
		.min(min10)		//交互比较后的最小的数据
	);										 
	switch switch11
	(
		//被比较交换的数输入
		.d0(max10),		//参与交互的第1个数
		.d1(min02),		//参与交互的第2个数
		//输出交互后的数据
		.max(max11),	//交互比较后的最大的数据
		.min(min11)		//交互比较后的最小的数据
	); 
	switch switch12
	(
		//被比较交换的数输入
		.d0(max11),		//参与交互的第1个数
		.d1(min03),		//参与交互的第2个数
		//输出交互后的数据
		.max(max12),	//交互比较后的最大的数据
		.min(min12)		//交互比较后的最小的数据
	);  
	switch switch13
	(
		//被比较交换的数输入
		.d0(max12),		//参与交互的第1个数
		.d1(min04),		//参与交互的第2个数
		//输出交互后的数据
		.max(max13),	//交互比较后的最大的数据
		.min(min13)		//交互比较后的最小的数据
	); 
	switch switch14
	(
		//被比较交换的数输入
		.d0(max13),		//参与交互的第1个数
		.d1(min05),		//参与交互的第2个数
		//输出交互后的数据
		.max(max14),	//交互比较后的最大的数据
		.min(min14)		//交互比较后的最小的数据
	); 
	switch switch15
	(
		//被比较交换的数输入
		.d0(max14),		//参与交互的第1个数
		.d1(min06),		//参与交互的第2个数
		//输出交互后的数据
		.max(max15),	//交互比较后的最大的数据
		.min(min15)		//交互比较后的最小的数据
	); 
	switch switch16
	(
		//被比较交换的数输入
		.d0(max15),		//参与交互的第1个数
		.d1(min07),		//参与交互的第2个数
		//输出交互后的数据
		.max(max16),	//交互比较后的最大的数据
		.min(min16)		//交互比较后的最小的数据
	);

	//第3次遍历/////////////
	wire [7:0] max20,max21,max22,max23,max24,max25;
	wire [7:0] min20,min21,min22,min23,min24,min25;
	switch switch20
	(
		//被比较交换的数输入
		.d0(min10),		//参与交互的第1个数
		.d1(min11),		//参与交互的第2个数
		//输出交互后的数据
		.max(max20),	//交互比较后的最大的数据
		.min(min20)		//交互比较后的最小的数据
	);
	switch switch21
	(
		//被比较交换的数输入
		.d0(max20),		//参与交互的第1个数
		.d1(min12),		//参与交互的第2个数
		//输出交互后的数据
		.max(max21),	//交互比较后的最大的数据
		.min(min21)		//交互比较后的最小的数据
	);	
	switch switch22
	(
		//被比较交换的数输入
		.d0(max21),		//参与交互的第1个数
		.d1(min13),		//参与交互的第2个数
		//输出交互后的数据
		.max(max22),	//交互比较后的最大的数据
		.min(min22)		//交互比较后的最小的数据
	);

	switch switch23
	(
		//被比较交换的数输入
		.d0(max22),		//参与交互的第1个数
		.d1(min14),		//参与交互的第2个数
		//输出交互后的数据
		.max(max23),	//交互比较后的最大的数据
		.min(min23)		//交互比较后的最小的数据
	);	
	switch switch24
	(
		//被比较交换的数输入
		.d0(max23),		//参与交互的第1个数
		.d1(min15),		//参与交互的第2个数
		//输出交互后的数据
		.max(max24),	//交互比较后的最大的数据
		.min(min24)		//交互比较后的最小的数据
	);	
	switch switch25
	(
		//被比较交换的数输入
		.d0(max24),		//参与交互的第1个数
		.d1(min16),		//参与交互的第2个数
		//输出交互后的数据
		.max(max25),	//交互比较后的最大的数据
		.min(min25)		//交互比较后的最小的数据
	);	

	//第4次遍历/////////////
	wire [7:0] max30,max31,max32,max33,max34;
	wire [7:0] min30,min31,min32,min33,min34;

	switch switch30
	(
		//被比较交换的数输入
		.d0(min20),		//参与交互的第1个数
		.d1(min21),		//参与交互的第2个数
		//输出交互后的数据
		.max(max30),	//交互比较后的最大的数据
		.min(min30)		//交互比较后的最小的数据
	);	
	switch switch31
	(
		//被比较交换的数输入
		.d0(max30),		//参与交互的第1个数
		.d1(min22),		//参与交互的第2个数
		//输出交互后的数据
		.max(max31),	//交互比较后的最大的数据
		.min(min31)		//交互比较后的最小的数据
	);
	switch switch32
	(
		//被比较交换的数输入
		.d0(max31),		//参与交互的第1个数
		.d1(min23),		//参与交互的第2个数
		//输出交互后的数据
		.max(max32),	//交互比较后的最大的数据
		.min(min32)		//交互比较后的最小的数据
	);	
	switch switch33
	(
		//被比较交换的数输入
		.d0(max32),		//参与交互的第1个数
		.d1(min24),		//参与交互的第2个数
		//输出交互后的数据
		.max(max33),	//交互比较后的最大的数据
		.min(min33)		//交互比较后的最小的数据
	);	
	switch switch34
	(
		//被比较交换的数输入
		.d0(max33),		//参与交互的第1个数
		.d1(min25),		//参与交互的第2个数
		//输出交互后的数据
		.max(max34),	//交互比较后的最大的数据
		.min(min34)		//交互比较后的最小的数据
	);

	//第5次遍历/////////////
	wire [7:0] max40,max41,max42,max43;
	wire [7:0] min40,min41,min42,min43;	
	switch switch40
	(
		//被比较交换的数输入
		.d0(min30),		//参与交互的第1个数
		.d1(min31),		//参与交互的第2个数
		//输出交互后的数据
		.max(max40),	//交互比较后的最大的数据
		.min(min40)		//交互比较后的最小的数据
	);

	switch switch41
	(
		//被比较交换的数输入
		.d0(max40),		//参与交互的第1个数
		.d1(min32),		//参与交互的第2个数
		//输出交互后的数据
		.max(max41),	//交互比较后的最大的数据
		.min(min41)		//交互比较后的最小的数据
	);
	switch switch42
	(
		//被比较交换的数输入
		.d0(max41),		//参与交互的第1个数
		.d1(min33),		//参与交互的第2个数
		//输出交互后的数据
		.max(max42),	//交互比较后的最大的数据
		.min(min42)		//交互比较后的最小的数据
	);
	switch switch43
	(
		//被比较交换的数输入
		.d0(max42),		//参与交互的第1个数
		.d1(min34),		//参与交互的第2个数
		//输出交互后的数据
		.max(max43),	//交互比较后的最大的数据
		.min(min43)		//交互比较后的最小的数据
	);

	assign oval[7:0] = max43[7:0];
endmodule