library verilog;
use verilog.vl_types.all;
entity vga565_sobel_tb is
end vga565_sobel_tb;
