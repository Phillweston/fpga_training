
module seven_tube_debug (
	source,
	probe);	

	output	[23:0]	source;
	input	[0:0]	probe;
endmodule
