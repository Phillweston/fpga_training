library verilog;
use verilog.vl_types.all;
entity crc_gen_tb is
end crc_gen_tb;
