module hour_flash ();
endmodule